 .GLOBAL vdd


 .TEMP 25.0
 .OPTION
 +    ARTIST=2
 +    INGOLD=2
 +    PARHIER=LOCAL
 +    PSF=2

 ** Library name: SPICE_Test
 ** Cell name: Diff_Amp_Basic
 ** View name: schematic
m1 net1 net2 net1 0 NMOS_VTL L=50e-9 W=90e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m2 net4 net5 net3 0 NMOS_VTL L=50e-9 W=90e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
m3 net5 net6 net2 0 NMOS_VTL L=50e-9 W=90e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
.END
